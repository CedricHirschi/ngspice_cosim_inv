** sch_path: /home/sem25f35/ngspice_cosim_inv/designs/comparator/comparator_tb.sch
**.subckt comparator_tb
x1 clk in_p in_n out2 out1 vss vdd comparator
Vdd vdd GND {vdd}
Vss vss GND {vss}
Vclk clk GND dc 0 ac 0 pulse({vss}, {vdd}, {0.9/f}, 1f, 1f, {0.1/f}, {1/f})
Vdiff in_p in_n pulse(2m, -2m, {0.75/f}, 1f, 1f, {1/f}, {2/f})
Vcm in_n GND {vdd/2}
E1 out1_dup GND VOL=' V(out1) '
E2 out2_dup GND VOL=' V(out2) '
XM5 out1_inv out1 vss vss sg13_lv_nmos w=1.5u l=0.13u ng=1 m=1
XM6 out1_inv out1 vdd vdd sg13_lv_pmos w=0.15u l=0.13u ng=1 m=1
XM7 out2_inv out2 vss vss sg13_lv_nmos w=1.5u l=0.13u ng=1 m=1
XM8 out2_inv out2 vdd vdd sg13_lv_pmos w=0.15u l=0.13u ng=1 m=1
XM1 out1_dup_inv out1_dup vss vss sg13_lv_nmos w=1.5u l=0.13u ng=1 m=1
XM2 out1_dup_inv out1_dup vdd vdd sg13_lv_pmos w=0.15u l=0.13u ng=1 m=1
XM3 out2_dup_inv out2_dup vss vss sg13_lv_nmos w=1.5u l=0.13u ng=1 m=1
XM4 out2_dup_inv out2_dup vdd vdd sg13_lv_pmos w=0.15u l=0.13u ng=1 m=1
**** begin user architecture code

.lib /foss/pdks/ihp-sg13g2/libs.tech/ngspice/models/cornerMOSlv.lib mos_tt
.include /foss/pdks/ihp-sg13g2/libs.ref/sg13g2_stdcell/spice/sg13g2_stdcell.spice




.param vss=0
.param vdd=1.5
.param f=100Meg

.tran 0.01n {4.5/f}


**** end user architecture code
**.ends

* expanding   symbol:  comparator.sym # of pins=7
** sym_path: /home/sem25f35/ngspice_cosim_inv/designs/comparator/comparator.sym
** sch_path: /home/sem25f35/ngspice_cosim_inv/designs/comparator/comparator.sch
.subckt comparator CLK IN1 IN2 OUT2 OUT1 VSS VDD
*.ipin CLK
*.ipin IN1
*.ipin IN2
*.opin OUT2
*.opin OUT1
*.ipin VSS
*.ipin VDD
XM1 net3 CLK VDD VDD sg13_lv_pmos w=2u l=0.13u ng=1 m=1
XM3 OUT1 OUT2 VDD VDD sg13_lv_pmos w=6u l=0.13u ng=3 m=1
XM4 OUT2 OUT1 VDD VDD sg13_lv_pmos w=6u l=0.13u ng=3 m=1
XM8 OUT1 OUT2 net3 VSS sg13_lv_nmos w=6u l=0.13u ng=3 m=1
XM9 net3 IN1 net1 VSS sg13_lv_nmos w=24u l=0.13u ng=12 m=1
XM11 net1 CLK VSS VSS sg13_lv_nmos w=24u l=0.26u ng=12 m=1
XM10 net2 IN2 net1 VSS sg13_lv_nmos w=24u l=0.13u ng=12 m=1
XM2 OUT1 CLK VDD VDD sg13_lv_pmos w=2u l=0.13u ng=1 m=1
XM5 net2 CLK VDD VDD sg13_lv_pmos w=2u l=0.13u ng=1 m=1
XM6 OUT2 CLK VDD VDD sg13_lv_pmos w=2u l=0.13u ng=1 m=1
XM7 OUT2 OUT1 net2 VSS sg13_lv_nmos w=6u l=0.13u ng=3 m=1
.ends

.GLOBAL GND
.end
